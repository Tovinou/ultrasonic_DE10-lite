-- watchdog_cpu_sys.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity watchdog_cpu_sys is
	port (
		button_export       : in    std_logic                     := '0';             --     button.export
		clk_clk             : in    std_logic                     := '0';             --        clk.clk
		hex_export          : out   std_logic_vector(6 downto 0);                     --        hex.export
		ledr_export         : out   std_logic_vector(7 downto 0);                     --       ledr.export
		pll_clk_clk         : out   std_logic;                                        --    pll_clk.clk
		reset_reset_n       : in    std_logic                     := '0';             --      reset.reset_n
		reset_out_reset_out : inout std_logic                     := '0';             --  reset_out.reset_out
		sdram_wire_addr     : out   std_logic_vector(12 downto 0);                    -- sdram_wire.addr
		sdram_wire_ba       : out   std_logic_vector(1 downto 0);                     --           .ba
		sdram_wire_cas_n    : out   std_logic;                                        --           .cas_n
		sdram_wire_cke      : out   std_logic;                                        --           .cke
		sdram_wire_cs_n     : out   std_logic;                                        --           .cs_n
		sdram_wire_dq       : inout std_logic_vector(15 downto 0) := (others => '0'); --           .dq
		sdram_wire_dqm      : out   std_logic_vector(1 downto 0);                     --           .dqm
		sdram_wire_ras_n    : out   std_logic;                                        --           .ras_n
		sdram_wire_we_n     : out   std_logic;                                        --           .we_n
		sw_export           : in    std_logic_vector(7 downto 0)  := (others => '0'); --         sw.export
		wdt_enable_export   : in    std_logic                     := '0'              -- wdt_enable.export
	);
end entity watchdog_cpu_sys;

architecture rtl of watchdog_cpu_sys is
	component watchdog_cpu_sys_CPU is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(27 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(27 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component watchdog_cpu_sys_CPU;

	component watchdog_cpu_sys_ENABLE is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic                     := 'X'              -- export
		);
	end component watchdog_cpu_sys_ENABLE;

	component watchdog_cpu_sys_LEDR is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component watchdog_cpu_sys_LEDR;

	component watchdog_cpu_sys_PIO_SWITCHES is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(7 downto 0)  := (others => 'X')  -- export
		);
	end component watchdog_cpu_sys_PIO_SWITCHES;

	component watchdog_cpu_sys_RAM is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(11 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component watchdog_cpu_sys_RAM;

	component watchdog_cpu_sys_SEVEN_SEG is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(6 downto 0)                      -- export
		);
	end component watchdog_cpu_sys_SEVEN_SEG;

	component TIMER_HW_IP is
		port (
			clk     : in  std_logic                     := 'X';             -- clk
			reset_n : in  std_logic                     := 'X';             -- reset_n
			cs_n    : in  std_logic                     := 'X';             -- chipselect_n
			addr    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n : in  std_logic                     := 'X';             -- write_n
			read_n  : in  std_logic                     := 'X';             -- read_n
			din     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dout    : out std_logic_vector(31 downto 0)                     -- readdata
		);
	end component TIMER_HW_IP;

	component WATCHDOG_TIMER_HW_IP is
		port (
			clk       : in    std_logic                     := 'X';             -- clk
			reset_n   : in    std_logic                     := 'X';             -- reset_n
			cs_n      : in    std_logic                     := 'X';             -- chipselect_n
			addr      : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n   : in    std_logic                     := 'X';             -- write_n
			read_n    : in    std_logic                     := 'X';             -- read_n
			din       : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dout      : out   std_logic_vector(31 downto 0);                    -- readdata
			reset_out : inout std_logic                     := 'X'              -- reset_out
		);
	end component WATCHDOG_TIMER_HW_IP;

	component watchdog_cpu_sys_altpll_0 is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			read               : in  std_logic                     := 'X';             -- read
			write              : in  std_logic                     := 'X';             -- write
			address            : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata           : out std_logic_vector(31 downto 0);                    -- readdata
			writedata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			c0                 : out std_logic;                                        -- clk
			c1                 : out std_logic;                                        -- clk
			scandone           : out std_logic;                                        -- export
			scandataout        : out std_logic;                                        -- export
			c2                 : out std_logic;                                        -- clk
			c3                 : out std_logic;                                        -- clk
			c4                 : out std_logic;                                        -- clk
			areset             : in  std_logic                     := 'X';             -- export
			locked             : out std_logic;                                        -- export
			phasedone          : out std_logic;                                        -- export
			phasecounterselect : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- export
			phaseupdown        : in  std_logic                     := 'X';             -- export
			phasestep          : in  std_logic                     := 'X';             -- export
			scanclk            : in  std_logic                     := 'X';             -- export
			scanclkena         : in  std_logic                     := 'X';             -- export
			scandata           : in  std_logic                     := 'X';             -- export
			configupdate       : in  std_logic                     := 'X'              -- export
		);
	end component watchdog_cpu_sys_altpll_0;

	component watchdog_cpu_sys_jtag_uart_0 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component watchdog_cpu_sys_jtag_uart_0;

	component watchdog_cpu_sys_sdram_controller is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(24 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component watchdog_cpu_sys_sdram_controller;

	component watchdog_cpu_sys_sysid_qsys_0 is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component watchdog_cpu_sys_sysid_qsys_0;

	component watchdog_cpu_sys_mm_interconnect_0 is
		port (
			altpll_0_c0_clk                                            : in  std_logic                     := 'X';             -- clk
			clk_0_clk_clk                                              : in  std_logic                     := 'X';             -- clk
			altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			CPU_reset_reset_bridge_in_reset_reset                      : in  std_logic                     := 'X';             -- reset
			CPU_data_master_address                                    : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			CPU_data_master_waitrequest                                : out std_logic;                                        -- waitrequest
			CPU_data_master_byteenable                                 : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			CPU_data_master_read                                       : in  std_logic                     := 'X';             -- read
			CPU_data_master_readdata                                   : out std_logic_vector(31 downto 0);                    -- readdata
			CPU_data_master_write                                      : in  std_logic                     := 'X';             -- write
			CPU_data_master_writedata                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			CPU_data_master_debugaccess                                : in  std_logic                     := 'X';             -- debugaccess
			CPU_instruction_master_address                             : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			CPU_instruction_master_waitrequest                         : out std_logic;                                        -- waitrequest
			CPU_instruction_master_read                                : in  std_logic                     := 'X';             -- read
			CPU_instruction_master_readdata                            : out std_logic_vector(31 downto 0);                    -- readdata
			altpll_0_pll_slave_address                                 : out std_logic_vector(1 downto 0);                     -- address
			altpll_0_pll_slave_write                                   : out std_logic;                                        -- write
			altpll_0_pll_slave_read                                    : out std_logic;                                        -- read
			altpll_0_pll_slave_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			altpll_0_pll_slave_writedata                               : out std_logic_vector(31 downto 0);                    -- writedata
			CPU_debug_mem_slave_address                                : out std_logic_vector(8 downto 0);                     -- address
			CPU_debug_mem_slave_write                                  : out std_logic;                                        -- write
			CPU_debug_mem_slave_read                                   : out std_logic;                                        -- read
			CPU_debug_mem_slave_readdata                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			CPU_debug_mem_slave_writedata                              : out std_logic_vector(31 downto 0);                    -- writedata
			CPU_debug_mem_slave_byteenable                             : out std_logic_vector(3 downto 0);                     -- byteenable
			CPU_debug_mem_slave_waitrequest                            : in  std_logic                     := 'X';             -- waitrequest
			CPU_debug_mem_slave_debugaccess                            : out std_logic;                                        -- debugaccess
			ENABLE_s1_address                                          : out std_logic_vector(1 downto 0);                     -- address
			ENABLE_s1_readdata                                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_0_avalon_jtag_slave_address                      : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_0_avalon_jtag_slave_write                        : out std_logic;                                        -- write
			jtag_uart_0_avalon_jtag_slave_read                         : out std_logic;                                        -- read
			jtag_uart_0_avalon_jtag_slave_readdata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_0_avalon_jtag_slave_writedata                    : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest                  : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect                   : out std_logic;                                        -- chipselect
			LEDR_s1_address                                            : out std_logic_vector(1 downto 0);                     -- address
			LEDR_s1_write                                              : out std_logic;                                        -- write
			LEDR_s1_readdata                                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			LEDR_s1_writedata                                          : out std_logic_vector(31 downto 0);                    -- writedata
			LEDR_s1_chipselect                                         : out std_logic;                                        -- chipselect
			PIO_BUTTON_s1_address                                      : out std_logic_vector(1 downto 0);                     -- address
			PIO_BUTTON_s1_readdata                                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			PIO_SWITCHES_s1_address                                    : out std_logic_vector(1 downto 0);                     -- address
			PIO_SWITCHES_s1_readdata                                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			RAM_s1_address                                             : out std_logic_vector(11 downto 0);                    -- address
			RAM_s1_write                                               : out std_logic;                                        -- write
			RAM_s1_readdata                                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			RAM_s1_writedata                                           : out std_logic_vector(31 downto 0);                    -- writedata
			RAM_s1_byteenable                                          : out std_logic_vector(3 downto 0);                     -- byteenable
			RAM_s1_chipselect                                          : out std_logic;                                        -- chipselect
			RAM_s1_clken                                               : out std_logic;                                        -- clken
			sdram_controller_s1_address                                : out std_logic_vector(24 downto 0);                    -- address
			sdram_controller_s1_write                                  : out std_logic;                                        -- write
			sdram_controller_s1_read                                   : out std_logic;                                        -- read
			sdram_controller_s1_readdata                               : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			sdram_controller_s1_writedata                              : out std_logic_vector(15 downto 0);                    -- writedata
			sdram_controller_s1_byteenable                             : out std_logic_vector(1 downto 0);                     -- byteenable
			sdram_controller_s1_readdatavalid                          : in  std_logic                     := 'X';             -- readdatavalid
			sdram_controller_s1_waitrequest                            : in  std_logic                     := 'X';             -- waitrequest
			sdram_controller_s1_chipselect                             : out std_logic;                                        -- chipselect
			SEVEN_SEG_s1_address                                       : out std_logic_vector(1 downto 0);                     -- address
			SEVEN_SEG_s1_write                                         : out std_logic;                                        -- write
			SEVEN_SEG_s1_readdata                                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			SEVEN_SEG_s1_writedata                                     : out std_logic_vector(31 downto 0);                    -- writedata
			SEVEN_SEG_s1_chipselect                                    : out std_logic;                                        -- chipselect
			sysid_qsys_0_control_slave_address                         : out std_logic_vector(0 downto 0);                     -- address
			sysid_qsys_0_control_slave_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			TIMER_HW_IP_0_avalon_slave_0_address                       : out std_logic_vector(1 downto 0);                     -- address
			TIMER_HW_IP_0_avalon_slave_0_write                         : out std_logic;                                        -- write
			TIMER_HW_IP_0_avalon_slave_0_read                          : out std_logic;                                        -- read
			TIMER_HW_IP_0_avalon_slave_0_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			TIMER_HW_IP_0_avalon_slave_0_writedata                     : out std_logic_vector(31 downto 0);                    -- writedata
			TIMER_HW_IP_0_avalon_slave_0_chipselect                    : out std_logic;                                        -- chipselect
			WATCHDOG_TIMER_HW_IP_0_avalon_slave_0_address              : out std_logic_vector(1 downto 0);                     -- address
			WATCHDOG_TIMER_HW_IP_0_avalon_slave_0_write                : out std_logic;                                        -- write
			WATCHDOG_TIMER_HW_IP_0_avalon_slave_0_read                 : out std_logic;                                        -- read
			WATCHDOG_TIMER_HW_IP_0_avalon_slave_0_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			WATCHDOG_TIMER_HW_IP_0_avalon_slave_0_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			WATCHDOG_TIMER_HW_IP_0_avalon_slave_0_chipselect           : out std_logic                                         -- chipselect
		);
	end component watchdog_cpu_sys_mm_interconnect_0;

	component watchdog_cpu_sys_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component watchdog_cpu_sys_irq_mapper;

	component watchdog_cpu_sys_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component watchdog_cpu_sys_rst_controller;

	component watchdog_cpu_sys_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component watchdog_cpu_sys_rst_controller_001;

	signal altpll_0_c0_clk                                                              : std_logic;                     -- altpll_0:c0 -> [CPU:clk, ENABLE:clk, LEDR:clk, PIO_BUTTON:clk, PIO_SWITCHES:clk, RAM:clk, SEVEN_SEG:clk, TIMER_HW_IP_0:clk, WATCHDOG_TIMER_HW_IP_0:clk, irq_mapper:clk, jtag_uart_0:clk, mm_interconnect_0:altpll_0_c0_clk, rst_controller:clk, sdram_controller:clk, sysid_qsys_0:clock]
	signal cpu_data_master_readdata                                                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:CPU_data_master_readdata -> CPU:d_readdata
	signal cpu_data_master_waitrequest                                                  : std_logic;                     -- mm_interconnect_0:CPU_data_master_waitrequest -> CPU:d_waitrequest
	signal cpu_data_master_debugaccess                                                  : std_logic;                     -- CPU:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:CPU_data_master_debugaccess
	signal cpu_data_master_address                                                      : std_logic_vector(27 downto 0); -- CPU:d_address -> mm_interconnect_0:CPU_data_master_address
	signal cpu_data_master_byteenable                                                   : std_logic_vector(3 downto 0);  -- CPU:d_byteenable -> mm_interconnect_0:CPU_data_master_byteenable
	signal cpu_data_master_read                                                         : std_logic;                     -- CPU:d_read -> mm_interconnect_0:CPU_data_master_read
	signal cpu_data_master_write                                                        : std_logic;                     -- CPU:d_write -> mm_interconnect_0:CPU_data_master_write
	signal cpu_data_master_writedata                                                    : std_logic_vector(31 downto 0); -- CPU:d_writedata -> mm_interconnect_0:CPU_data_master_writedata
	signal cpu_instruction_master_readdata                                              : std_logic_vector(31 downto 0); -- mm_interconnect_0:CPU_instruction_master_readdata -> CPU:i_readdata
	signal cpu_instruction_master_waitrequest                                           : std_logic;                     -- mm_interconnect_0:CPU_instruction_master_waitrequest -> CPU:i_waitrequest
	signal cpu_instruction_master_address                                               : std_logic_vector(27 downto 0); -- CPU:i_address -> mm_interconnect_0:CPU_instruction_master_address
	signal cpu_instruction_master_read                                                  : std_logic;                     -- CPU:i_read -> mm_interconnect_0:CPU_instruction_master_read
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect                   : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata                     : std_logic_vector(31 downto 0); -- jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest                  : std_logic;                     -- jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address                      : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read                         : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write                        : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	signal mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_chipselect                    : std_logic;                     -- mm_interconnect_0:TIMER_HW_IP_0_avalon_slave_0_chipselect -> mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_chipselect:in
	signal mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_readdata                      : std_logic_vector(31 downto 0); -- TIMER_HW_IP_0:dout -> mm_interconnect_0:TIMER_HW_IP_0_avalon_slave_0_readdata
	signal mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_address                       : std_logic_vector(1 downto 0);  -- mm_interconnect_0:TIMER_HW_IP_0_avalon_slave_0_address -> TIMER_HW_IP_0:addr
	signal mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_read                          : std_logic;                     -- mm_interconnect_0:TIMER_HW_IP_0_avalon_slave_0_read -> mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_read:in
	signal mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_write                         : std_logic;                     -- mm_interconnect_0:TIMER_HW_IP_0_avalon_slave_0_write -> mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_write:in
	signal mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_writedata                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:TIMER_HW_IP_0_avalon_slave_0_writedata -> TIMER_HW_IP_0:din
	signal mm_interconnect_0_watchdog_timer_hw_ip_0_avalon_slave_0_chipselect           : std_logic;                     -- mm_interconnect_0:WATCHDOG_TIMER_HW_IP_0_avalon_slave_0_chipselect -> mm_interconnect_0_watchdog_timer_hw_ip_0_avalon_slave_0_chipselect:in
	signal mm_interconnect_0_watchdog_timer_hw_ip_0_avalon_slave_0_readdata             : std_logic_vector(31 downto 0); -- WATCHDOG_TIMER_HW_IP_0:dout -> mm_interconnect_0:WATCHDOG_TIMER_HW_IP_0_avalon_slave_0_readdata
	signal mm_interconnect_0_watchdog_timer_hw_ip_0_avalon_slave_0_address              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:WATCHDOG_TIMER_HW_IP_0_avalon_slave_0_address -> WATCHDOG_TIMER_HW_IP_0:addr
	signal mm_interconnect_0_watchdog_timer_hw_ip_0_avalon_slave_0_read                 : std_logic;                     -- mm_interconnect_0:WATCHDOG_TIMER_HW_IP_0_avalon_slave_0_read -> mm_interconnect_0_watchdog_timer_hw_ip_0_avalon_slave_0_read:in
	signal mm_interconnect_0_watchdog_timer_hw_ip_0_avalon_slave_0_write                : std_logic;                     -- mm_interconnect_0:WATCHDOG_TIMER_HW_IP_0_avalon_slave_0_write -> mm_interconnect_0_watchdog_timer_hw_ip_0_avalon_slave_0_write:in
	signal mm_interconnect_0_watchdog_timer_hw_ip_0_avalon_slave_0_writedata            : std_logic_vector(31 downto 0); -- mm_interconnect_0:WATCHDOG_TIMER_HW_IP_0_avalon_slave_0_writedata -> WATCHDOG_TIMER_HW_IP_0:din
	signal mm_interconnect_0_sysid_qsys_0_control_slave_readdata                        : std_logic_vector(31 downto 0); -- sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	signal mm_interconnect_0_sysid_qsys_0_control_slave_address                         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	signal mm_interconnect_0_cpu_debug_mem_slave_readdata                               : std_logic_vector(31 downto 0); -- CPU:debug_mem_slave_readdata -> mm_interconnect_0:CPU_debug_mem_slave_readdata
	signal mm_interconnect_0_cpu_debug_mem_slave_waitrequest                            : std_logic;                     -- CPU:debug_mem_slave_waitrequest -> mm_interconnect_0:CPU_debug_mem_slave_waitrequest
	signal mm_interconnect_0_cpu_debug_mem_slave_debugaccess                            : std_logic;                     -- mm_interconnect_0:CPU_debug_mem_slave_debugaccess -> CPU:debug_mem_slave_debugaccess
	signal mm_interconnect_0_cpu_debug_mem_slave_address                                : std_logic_vector(8 downto 0);  -- mm_interconnect_0:CPU_debug_mem_slave_address -> CPU:debug_mem_slave_address
	signal mm_interconnect_0_cpu_debug_mem_slave_read                                   : std_logic;                     -- mm_interconnect_0:CPU_debug_mem_slave_read -> CPU:debug_mem_slave_read
	signal mm_interconnect_0_cpu_debug_mem_slave_byteenable                             : std_logic_vector(3 downto 0);  -- mm_interconnect_0:CPU_debug_mem_slave_byteenable -> CPU:debug_mem_slave_byteenable
	signal mm_interconnect_0_cpu_debug_mem_slave_write                                  : std_logic;                     -- mm_interconnect_0:CPU_debug_mem_slave_write -> CPU:debug_mem_slave_write
	signal mm_interconnect_0_cpu_debug_mem_slave_writedata                              : std_logic_vector(31 downto 0); -- mm_interconnect_0:CPU_debug_mem_slave_writedata -> CPU:debug_mem_slave_writedata
	signal mm_interconnect_0_altpll_0_pll_slave_readdata                                : std_logic_vector(31 downto 0); -- altpll_0:readdata -> mm_interconnect_0:altpll_0_pll_slave_readdata
	signal mm_interconnect_0_altpll_0_pll_slave_address                                 : std_logic_vector(1 downto 0);  -- mm_interconnect_0:altpll_0_pll_slave_address -> altpll_0:address
	signal mm_interconnect_0_altpll_0_pll_slave_read                                    : std_logic;                     -- mm_interconnect_0:altpll_0_pll_slave_read -> altpll_0:read
	signal mm_interconnect_0_altpll_0_pll_slave_write                                   : std_logic;                     -- mm_interconnect_0:altpll_0_pll_slave_write -> altpll_0:write
	signal mm_interconnect_0_altpll_0_pll_slave_writedata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:altpll_0_pll_slave_writedata -> altpll_0:writedata
	signal mm_interconnect_0_ram_s1_chipselect                                          : std_logic;                     -- mm_interconnect_0:RAM_s1_chipselect -> RAM:chipselect
	signal mm_interconnect_0_ram_s1_readdata                                            : std_logic_vector(31 downto 0); -- RAM:readdata -> mm_interconnect_0:RAM_s1_readdata
	signal mm_interconnect_0_ram_s1_address                                             : std_logic_vector(11 downto 0); -- mm_interconnect_0:RAM_s1_address -> RAM:address
	signal mm_interconnect_0_ram_s1_byteenable                                          : std_logic_vector(3 downto 0);  -- mm_interconnect_0:RAM_s1_byteenable -> RAM:byteenable
	signal mm_interconnect_0_ram_s1_write                                               : std_logic;                     -- mm_interconnect_0:RAM_s1_write -> RAM:write
	signal mm_interconnect_0_ram_s1_writedata                                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:RAM_s1_writedata -> RAM:writedata
	signal mm_interconnect_0_ram_s1_clken                                               : std_logic;                     -- mm_interconnect_0:RAM_s1_clken -> RAM:clken
	signal mm_interconnect_0_pio_switches_s1_readdata                                   : std_logic_vector(31 downto 0); -- PIO_SWITCHES:readdata -> mm_interconnect_0:PIO_SWITCHES_s1_readdata
	signal mm_interconnect_0_pio_switches_s1_address                                    : std_logic_vector(1 downto 0);  -- mm_interconnect_0:PIO_SWITCHES_s1_address -> PIO_SWITCHES:address
	signal mm_interconnect_0_pio_button_s1_readdata                                     : std_logic_vector(31 downto 0); -- PIO_BUTTON:readdata -> mm_interconnect_0:PIO_BUTTON_s1_readdata
	signal mm_interconnect_0_pio_button_s1_address                                      : std_logic_vector(1 downto 0);  -- mm_interconnect_0:PIO_BUTTON_s1_address -> PIO_BUTTON:address
	signal mm_interconnect_0_ledr_s1_chipselect                                         : std_logic;                     -- mm_interconnect_0:LEDR_s1_chipselect -> LEDR:chipselect
	signal mm_interconnect_0_ledr_s1_readdata                                           : std_logic_vector(31 downto 0); -- LEDR:readdata -> mm_interconnect_0:LEDR_s1_readdata
	signal mm_interconnect_0_ledr_s1_address                                            : std_logic_vector(1 downto 0);  -- mm_interconnect_0:LEDR_s1_address -> LEDR:address
	signal mm_interconnect_0_ledr_s1_write                                              : std_logic;                     -- mm_interconnect_0:LEDR_s1_write -> mm_interconnect_0_ledr_s1_write:in
	signal mm_interconnect_0_ledr_s1_writedata                                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:LEDR_s1_writedata -> LEDR:writedata
	signal mm_interconnect_0_seven_seg_s1_chipselect                                    : std_logic;                     -- mm_interconnect_0:SEVEN_SEG_s1_chipselect -> SEVEN_SEG:chipselect
	signal mm_interconnect_0_seven_seg_s1_readdata                                      : std_logic_vector(31 downto 0); -- SEVEN_SEG:readdata -> mm_interconnect_0:SEVEN_SEG_s1_readdata
	signal mm_interconnect_0_seven_seg_s1_address                                       : std_logic_vector(1 downto 0);  -- mm_interconnect_0:SEVEN_SEG_s1_address -> SEVEN_SEG:address
	signal mm_interconnect_0_seven_seg_s1_write                                         : std_logic;                     -- mm_interconnect_0:SEVEN_SEG_s1_write -> mm_interconnect_0_seven_seg_s1_write:in
	signal mm_interconnect_0_seven_seg_s1_writedata                                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:SEVEN_SEG_s1_writedata -> SEVEN_SEG:writedata
	signal mm_interconnect_0_enable_s1_readdata                                         : std_logic_vector(31 downto 0); -- ENABLE:readdata -> mm_interconnect_0:ENABLE_s1_readdata
	signal mm_interconnect_0_enable_s1_address                                          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:ENABLE_s1_address -> ENABLE:address
	signal mm_interconnect_0_sdram_controller_s1_chipselect                             : std_logic;                     -- mm_interconnect_0:sdram_controller_s1_chipselect -> sdram_controller:az_cs
	signal mm_interconnect_0_sdram_controller_s1_readdata                               : std_logic_vector(15 downto 0); -- sdram_controller:za_data -> mm_interconnect_0:sdram_controller_s1_readdata
	signal mm_interconnect_0_sdram_controller_s1_waitrequest                            : std_logic;                     -- sdram_controller:za_waitrequest -> mm_interconnect_0:sdram_controller_s1_waitrequest
	signal mm_interconnect_0_sdram_controller_s1_address                                : std_logic_vector(24 downto 0); -- mm_interconnect_0:sdram_controller_s1_address -> sdram_controller:az_addr
	signal mm_interconnect_0_sdram_controller_s1_read                                   : std_logic;                     -- mm_interconnect_0:sdram_controller_s1_read -> mm_interconnect_0_sdram_controller_s1_read:in
	signal mm_interconnect_0_sdram_controller_s1_byteenable                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:sdram_controller_s1_byteenable -> mm_interconnect_0_sdram_controller_s1_byteenable:in
	signal mm_interconnect_0_sdram_controller_s1_readdatavalid                          : std_logic;                     -- sdram_controller:za_valid -> mm_interconnect_0:sdram_controller_s1_readdatavalid
	signal mm_interconnect_0_sdram_controller_s1_write                                  : std_logic;                     -- mm_interconnect_0:sdram_controller_s1_write -> mm_interconnect_0_sdram_controller_s1_write:in
	signal mm_interconnect_0_sdram_controller_s1_writedata                              : std_logic_vector(15 downto 0); -- mm_interconnect_0:sdram_controller_s1_writedata -> sdram_controller:az_data
	signal irq_mapper_receiver0_irq                                                     : std_logic;                     -- jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	signal cpu_irq_irq                                                                  : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> CPU:irq
	signal rst_controller_reset_out_reset                                               : std_logic;                     -- rst_controller:reset_out -> [RAM:reset, irq_mapper:reset, mm_interconnect_0:CPU_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                                           : std_logic;                     -- rst_controller:reset_req -> [CPU:reset_req, RAM:reset_req, rst_translator:reset_req_in]
	signal cpu_debug_reset_request_reset                                                : std_logic;                     -- CPU:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	signal rst_controller_001_reset_out_reset                                           : std_logic;                     -- rst_controller_001:reset_out -> [altpll_0:reset, mm_interconnect_0:altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset]
	signal reset_reset_n_ports_inv                                                      : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0]
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv               : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:inv -> jtag_uart_0:av_read_n
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv              : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:inv -> jtag_uart_0:av_write_n
	signal mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_chipselect_ports_inv          : std_logic;                     -- mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_chipselect:inv -> TIMER_HW_IP_0:cs_n
	signal mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_read_ports_inv                : std_logic;                     -- mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_read:inv -> TIMER_HW_IP_0:read_n
	signal mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_write_ports_inv               : std_logic;                     -- mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_write:inv -> TIMER_HW_IP_0:write_n
	signal mm_interconnect_0_watchdog_timer_hw_ip_0_avalon_slave_0_chipselect_ports_inv : std_logic;                     -- mm_interconnect_0_watchdog_timer_hw_ip_0_avalon_slave_0_chipselect:inv -> WATCHDOG_TIMER_HW_IP_0:cs_n
	signal mm_interconnect_0_watchdog_timer_hw_ip_0_avalon_slave_0_read_ports_inv       : std_logic;                     -- mm_interconnect_0_watchdog_timer_hw_ip_0_avalon_slave_0_read:inv -> WATCHDOG_TIMER_HW_IP_0:read_n
	signal mm_interconnect_0_watchdog_timer_hw_ip_0_avalon_slave_0_write_ports_inv      : std_logic;                     -- mm_interconnect_0_watchdog_timer_hw_ip_0_avalon_slave_0_write:inv -> WATCHDOG_TIMER_HW_IP_0:write_n
	signal mm_interconnect_0_ledr_s1_write_ports_inv                                    : std_logic;                     -- mm_interconnect_0_ledr_s1_write:inv -> LEDR:write_n
	signal mm_interconnect_0_seven_seg_s1_write_ports_inv                               : std_logic;                     -- mm_interconnect_0_seven_seg_s1_write:inv -> SEVEN_SEG:write_n
	signal mm_interconnect_0_sdram_controller_s1_read_ports_inv                         : std_logic;                     -- mm_interconnect_0_sdram_controller_s1_read:inv -> sdram_controller:az_rd_n
	signal mm_interconnect_0_sdram_controller_s1_byteenable_ports_inv                   : std_logic_vector(1 downto 0);  -- mm_interconnect_0_sdram_controller_s1_byteenable:inv -> sdram_controller:az_be_n
	signal mm_interconnect_0_sdram_controller_s1_write_ports_inv                        : std_logic;                     -- mm_interconnect_0_sdram_controller_s1_write:inv -> sdram_controller:az_wr_n
	signal rst_controller_reset_out_reset_ports_inv                                     : std_logic;                     -- rst_controller_reset_out_reset:inv -> [CPU:reset_n, ENABLE:reset_n, LEDR:reset_n, PIO_BUTTON:reset_n, PIO_SWITCHES:reset_n, SEVEN_SEG:reset_n, TIMER_HW_IP_0:reset_n, WATCHDOG_TIMER_HW_IP_0:reset_n, jtag_uart_0:rst_n, sdram_controller:reset_n, sysid_qsys_0:reset_n]

begin

	cpu : component watchdog_cpu_sys_CPU
		port map (
			clk                                 => altpll_0_c0_clk,                                   --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,          --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                --                          .reset_req
			d_address                           => cpu_data_master_address,                           --               data_master.address
			d_byteenable                        => cpu_data_master_byteenable,                        --                          .byteenable
			d_read                              => cpu_data_master_read,                              --                          .read
			d_readdata                          => cpu_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => cpu_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => cpu_data_master_write,                             --                          .write
			d_writedata                         => cpu_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => cpu_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => cpu_instruction_master_address,                    --        instruction_master.address
			i_read                              => cpu_instruction_master_read,                       --                          .read
			i_readdata                          => cpu_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => cpu_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => cpu_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => cpu_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_cpu_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_cpu_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_cpu_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_cpu_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_cpu_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_cpu_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_cpu_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_cpu_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                               -- custom_instruction_master.readra
		);

	enable : component watchdog_cpu_sys_ENABLE
		port map (
			clk      => altpll_0_c0_clk,                          --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_enable_s1_address,      --                  s1.address
			readdata => mm_interconnect_0_enable_s1_readdata,     --                    .readdata
			in_port  => wdt_enable_export                         -- external_connection.export
		);

	ledr : component watchdog_cpu_sys_LEDR
		port map (
			clk        => altpll_0_c0_clk,                           --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_0_ledr_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_ledr_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_ledr_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_ledr_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_ledr_s1_readdata,        --                    .readdata
			out_port   => ledr_export                                -- external_connection.export
		);

	pio_button : component watchdog_cpu_sys_ENABLE
		port map (
			clk      => altpll_0_c0_clk,                          --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_pio_button_s1_address,  --                  s1.address
			readdata => mm_interconnect_0_pio_button_s1_readdata, --                    .readdata
			in_port  => button_export                             -- external_connection.export
		);

	pio_switches : component watchdog_cpu_sys_PIO_SWITCHES
		port map (
			clk      => altpll_0_c0_clk,                            --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address  => mm_interconnect_0_pio_switches_s1_address,  --                  s1.address
			readdata => mm_interconnect_0_pio_switches_s1_readdata, --                    .readdata
			in_port  => sw_export                                   -- external_connection.export
		);

	ram : component watchdog_cpu_sys_RAM
		port map (
			clk        => altpll_0_c0_clk,                     --   clk1.clk
			address    => mm_interconnect_0_ram_s1_address,    --     s1.address
			clken      => mm_interconnect_0_ram_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_ram_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_ram_s1_write,      --       .write
			readdata   => mm_interconnect_0_ram_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_ram_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_ram_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,      -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,  --       .reset_req
			freeze     => '0'                                  -- (terminated)
		);

	seven_seg : component watchdog_cpu_sys_SEVEN_SEG
		port map (
			clk        => altpll_0_c0_clk,                                --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,       --               reset.reset_n
			address    => mm_interconnect_0_seven_seg_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_seven_seg_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_seven_seg_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_seven_seg_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_seven_seg_s1_readdata,        --                    .readdata
			out_port   => hex_export                                      -- external_connection.export
		);

	timer_hw_ip_0 : component TIMER_HW_IP
		port map (
			clk     => altpll_0_c0_clk,                                                     --          clock.clk
			reset_n => rst_controller_reset_out_reset_ports_inv,                            --          reset.reset_n
			cs_n    => mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_chipselect_ports_inv, -- avalon_slave_0.chipselect_n
			addr    => mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_address,              --               .address
			write_n => mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_write_ports_inv,      --               .write_n
			read_n  => mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_read_ports_inv,       --               .read_n
			din     => mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_writedata,            --               .writedata
			dout    => mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_readdata              --               .readdata
		);

	watchdog_timer_hw_ip_0 : component WATCHDOG_TIMER_HW_IP
		port map (
			clk       => altpll_0_c0_clk,                                                              --          clock.clk
			reset_n   => rst_controller_reset_out_reset_ports_inv,                                     --          reset.reset_n
			cs_n      => mm_interconnect_0_watchdog_timer_hw_ip_0_avalon_slave_0_chipselect_ports_inv, -- avalon_slave_0.chipselect_n
			addr      => mm_interconnect_0_watchdog_timer_hw_ip_0_avalon_slave_0_address,              --               .address
			write_n   => mm_interconnect_0_watchdog_timer_hw_ip_0_avalon_slave_0_write_ports_inv,      --               .write_n
			read_n    => mm_interconnect_0_watchdog_timer_hw_ip_0_avalon_slave_0_read_ports_inv,       --               .read_n
			din       => mm_interconnect_0_watchdog_timer_hw_ip_0_avalon_slave_0_writedata,            --               .writedata
			dout      => mm_interconnect_0_watchdog_timer_hw_ip_0_avalon_slave_0_readdata,             --               .readdata
			reset_out => reset_out_reset_out                                                           --    conduit_end.reset_out
		);

	altpll_0 : component watchdog_cpu_sys_altpll_0
		port map (
			clk                => clk_clk,                                        --       inclk_interface.clk
			reset              => rst_controller_001_reset_out_reset,             -- inclk_interface_reset.reset
			read               => mm_interconnect_0_altpll_0_pll_slave_read,      --             pll_slave.read
			write              => mm_interconnect_0_altpll_0_pll_slave_write,     --                      .write
			address            => mm_interconnect_0_altpll_0_pll_slave_address,   --                      .address
			readdata           => mm_interconnect_0_altpll_0_pll_slave_readdata,  --                      .readdata
			writedata          => mm_interconnect_0_altpll_0_pll_slave_writedata, --                      .writedata
			c0                 => altpll_0_c0_clk,                                --                    c0.clk
			c1                 => pll_clk_clk,                                    --                    c1.clk
			scandone           => open,                                           --           (terminated)
			scandataout        => open,                                           --           (terminated)
			c2                 => open,                                           --           (terminated)
			c3                 => open,                                           --           (terminated)
			c4                 => open,                                           --           (terminated)
			areset             => '0',                                            --           (terminated)
			locked             => open,                                           --           (terminated)
			phasedone          => open,                                           --           (terminated)
			phasecounterselect => "000",                                          --           (terminated)
			phaseupdown        => '0',                                            --           (terminated)
			phasestep          => '0',                                            --           (terminated)
			scanclk            => '0',                                            --           (terminated)
			scanclkena         => '0',                                            --           (terminated)
			scandata           => '0',                                            --           (terminated)
			configupdate       => '0'                                             --           (terminated)
		);

	jtag_uart_0 : component watchdog_cpu_sys_jtag_uart_0
		port map (
			clk            => altpll_0_c0_clk,                                                 --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                        --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                         --               irq.irq
		);

	sdram_controller : component watchdog_cpu_sys_sdram_controller
		port map (
			clk            => altpll_0_c0_clk,                                            --   clk.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,                   -- reset.reset_n
			az_addr        => mm_interconnect_0_sdram_controller_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_sdram_controller_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_sdram_controller_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_sdram_controller_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_sdram_controller_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_sdram_controller_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_sdram_controller_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_sdram_controller_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_sdram_controller_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_wire_addr,                                            --  wire.export
			zs_ba          => sdram_wire_ba,                                              --      .export
			zs_cas_n       => sdram_wire_cas_n,                                           --      .export
			zs_cke         => sdram_wire_cke,                                             --      .export
			zs_cs_n        => sdram_wire_cs_n,                                            --      .export
			zs_dq          => sdram_wire_dq,                                              --      .export
			zs_dqm         => sdram_wire_dqm,                                             --      .export
			zs_ras_n       => sdram_wire_ras_n,                                           --      .export
			zs_we_n        => sdram_wire_we_n                                             --      .export
		);

	sysid_qsys_0 : component watchdog_cpu_sys_sysid_qsys_0
		port map (
			clock    => altpll_0_c0_clk,                                         --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,                --         reset.reset_n
			readdata => mm_interconnect_0_sysid_qsys_0_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_qsys_0_control_slave_address(0)  --              .address
		);

	mm_interconnect_0 : component watchdog_cpu_sys_mm_interconnect_0
		port map (
			altpll_0_c0_clk                                            => altpll_0_c0_clk,                                                    --                                          altpll_0_c0.clk
			clk_0_clk_clk                                              => clk_clk,                                                            --                                            clk_0_clk.clk
			altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset => rst_controller_001_reset_out_reset,                                 -- altpll_0_inclk_interface_reset_reset_bridge_in_reset.reset
			CPU_reset_reset_bridge_in_reset_reset                      => rst_controller_reset_out_reset,                                     --                      CPU_reset_reset_bridge_in_reset.reset
			CPU_data_master_address                                    => cpu_data_master_address,                                            --                                      CPU_data_master.address
			CPU_data_master_waitrequest                                => cpu_data_master_waitrequest,                                        --                                                     .waitrequest
			CPU_data_master_byteenable                                 => cpu_data_master_byteenable,                                         --                                                     .byteenable
			CPU_data_master_read                                       => cpu_data_master_read,                                               --                                                     .read
			CPU_data_master_readdata                                   => cpu_data_master_readdata,                                           --                                                     .readdata
			CPU_data_master_write                                      => cpu_data_master_write,                                              --                                                     .write
			CPU_data_master_writedata                                  => cpu_data_master_writedata,                                          --                                                     .writedata
			CPU_data_master_debugaccess                                => cpu_data_master_debugaccess,                                        --                                                     .debugaccess
			CPU_instruction_master_address                             => cpu_instruction_master_address,                                     --                               CPU_instruction_master.address
			CPU_instruction_master_waitrequest                         => cpu_instruction_master_waitrequest,                                 --                                                     .waitrequest
			CPU_instruction_master_read                                => cpu_instruction_master_read,                                        --                                                     .read
			CPU_instruction_master_readdata                            => cpu_instruction_master_readdata,                                    --                                                     .readdata
			altpll_0_pll_slave_address                                 => mm_interconnect_0_altpll_0_pll_slave_address,                       --                                   altpll_0_pll_slave.address
			altpll_0_pll_slave_write                                   => mm_interconnect_0_altpll_0_pll_slave_write,                         --                                                     .write
			altpll_0_pll_slave_read                                    => mm_interconnect_0_altpll_0_pll_slave_read,                          --                                                     .read
			altpll_0_pll_slave_readdata                                => mm_interconnect_0_altpll_0_pll_slave_readdata,                      --                                                     .readdata
			altpll_0_pll_slave_writedata                               => mm_interconnect_0_altpll_0_pll_slave_writedata,                     --                                                     .writedata
			CPU_debug_mem_slave_address                                => mm_interconnect_0_cpu_debug_mem_slave_address,                      --                                  CPU_debug_mem_slave.address
			CPU_debug_mem_slave_write                                  => mm_interconnect_0_cpu_debug_mem_slave_write,                        --                                                     .write
			CPU_debug_mem_slave_read                                   => mm_interconnect_0_cpu_debug_mem_slave_read,                         --                                                     .read
			CPU_debug_mem_slave_readdata                               => mm_interconnect_0_cpu_debug_mem_slave_readdata,                     --                                                     .readdata
			CPU_debug_mem_slave_writedata                              => mm_interconnect_0_cpu_debug_mem_slave_writedata,                    --                                                     .writedata
			CPU_debug_mem_slave_byteenable                             => mm_interconnect_0_cpu_debug_mem_slave_byteenable,                   --                                                     .byteenable
			CPU_debug_mem_slave_waitrequest                            => mm_interconnect_0_cpu_debug_mem_slave_waitrequest,                  --                                                     .waitrequest
			CPU_debug_mem_slave_debugaccess                            => mm_interconnect_0_cpu_debug_mem_slave_debugaccess,                  --                                                     .debugaccess
			ENABLE_s1_address                                          => mm_interconnect_0_enable_s1_address,                                --                                            ENABLE_s1.address
			ENABLE_s1_readdata                                         => mm_interconnect_0_enable_s1_readdata,                               --                                                     .readdata
			jtag_uart_0_avalon_jtag_slave_address                      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address,            --                        jtag_uart_0_avalon_jtag_slave.address
			jtag_uart_0_avalon_jtag_slave_write                        => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write,              --                                                     .write
			jtag_uart_0_avalon_jtag_slave_read                         => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read,               --                                                     .read
			jtag_uart_0_avalon_jtag_slave_readdata                     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,           --                                                     .readdata
			jtag_uart_0_avalon_jtag_slave_writedata                    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,          --                                                     .writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest                  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,        --                                                     .waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect                   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,         --                                                     .chipselect
			LEDR_s1_address                                            => mm_interconnect_0_ledr_s1_address,                                  --                                              LEDR_s1.address
			LEDR_s1_write                                              => mm_interconnect_0_ledr_s1_write,                                    --                                                     .write
			LEDR_s1_readdata                                           => mm_interconnect_0_ledr_s1_readdata,                                 --                                                     .readdata
			LEDR_s1_writedata                                          => mm_interconnect_0_ledr_s1_writedata,                                --                                                     .writedata
			LEDR_s1_chipselect                                         => mm_interconnect_0_ledr_s1_chipselect,                               --                                                     .chipselect
			PIO_BUTTON_s1_address                                      => mm_interconnect_0_pio_button_s1_address,                            --                                        PIO_BUTTON_s1.address
			PIO_BUTTON_s1_readdata                                     => mm_interconnect_0_pio_button_s1_readdata,                           --                                                     .readdata
			PIO_SWITCHES_s1_address                                    => mm_interconnect_0_pio_switches_s1_address,                          --                                      PIO_SWITCHES_s1.address
			PIO_SWITCHES_s1_readdata                                   => mm_interconnect_0_pio_switches_s1_readdata,                         --                                                     .readdata
			RAM_s1_address                                             => mm_interconnect_0_ram_s1_address,                                   --                                               RAM_s1.address
			RAM_s1_write                                               => mm_interconnect_0_ram_s1_write,                                     --                                                     .write
			RAM_s1_readdata                                            => mm_interconnect_0_ram_s1_readdata,                                  --                                                     .readdata
			RAM_s1_writedata                                           => mm_interconnect_0_ram_s1_writedata,                                 --                                                     .writedata
			RAM_s1_byteenable                                          => mm_interconnect_0_ram_s1_byteenable,                                --                                                     .byteenable
			RAM_s1_chipselect                                          => mm_interconnect_0_ram_s1_chipselect,                                --                                                     .chipselect
			RAM_s1_clken                                               => mm_interconnect_0_ram_s1_clken,                                     --                                                     .clken
			sdram_controller_s1_address                                => mm_interconnect_0_sdram_controller_s1_address,                      --                                  sdram_controller_s1.address
			sdram_controller_s1_write                                  => mm_interconnect_0_sdram_controller_s1_write,                        --                                                     .write
			sdram_controller_s1_read                                   => mm_interconnect_0_sdram_controller_s1_read,                         --                                                     .read
			sdram_controller_s1_readdata                               => mm_interconnect_0_sdram_controller_s1_readdata,                     --                                                     .readdata
			sdram_controller_s1_writedata                              => mm_interconnect_0_sdram_controller_s1_writedata,                    --                                                     .writedata
			sdram_controller_s1_byteenable                             => mm_interconnect_0_sdram_controller_s1_byteenable,                   --                                                     .byteenable
			sdram_controller_s1_readdatavalid                          => mm_interconnect_0_sdram_controller_s1_readdatavalid,                --                                                     .readdatavalid
			sdram_controller_s1_waitrequest                            => mm_interconnect_0_sdram_controller_s1_waitrequest,                  --                                                     .waitrequest
			sdram_controller_s1_chipselect                             => mm_interconnect_0_sdram_controller_s1_chipselect,                   --                                                     .chipselect
			SEVEN_SEG_s1_address                                       => mm_interconnect_0_seven_seg_s1_address,                             --                                         SEVEN_SEG_s1.address
			SEVEN_SEG_s1_write                                         => mm_interconnect_0_seven_seg_s1_write,                               --                                                     .write
			SEVEN_SEG_s1_readdata                                      => mm_interconnect_0_seven_seg_s1_readdata,                            --                                                     .readdata
			SEVEN_SEG_s1_writedata                                     => mm_interconnect_0_seven_seg_s1_writedata,                           --                                                     .writedata
			SEVEN_SEG_s1_chipselect                                    => mm_interconnect_0_seven_seg_s1_chipselect,                          --                                                     .chipselect
			sysid_qsys_0_control_slave_address                         => mm_interconnect_0_sysid_qsys_0_control_slave_address,               --                           sysid_qsys_0_control_slave.address
			sysid_qsys_0_control_slave_readdata                        => mm_interconnect_0_sysid_qsys_0_control_slave_readdata,              --                                                     .readdata
			TIMER_HW_IP_0_avalon_slave_0_address                       => mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_address,             --                         TIMER_HW_IP_0_avalon_slave_0.address
			TIMER_HW_IP_0_avalon_slave_0_write                         => mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_write,               --                                                     .write
			TIMER_HW_IP_0_avalon_slave_0_read                          => mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_read,                --                                                     .read
			TIMER_HW_IP_0_avalon_slave_0_readdata                      => mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_readdata,            --                                                     .readdata
			TIMER_HW_IP_0_avalon_slave_0_writedata                     => mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_writedata,           --                                                     .writedata
			TIMER_HW_IP_0_avalon_slave_0_chipselect                    => mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_chipselect,          --                                                     .chipselect
			WATCHDOG_TIMER_HW_IP_0_avalon_slave_0_address              => mm_interconnect_0_watchdog_timer_hw_ip_0_avalon_slave_0_address,    --                WATCHDOG_TIMER_HW_IP_0_avalon_slave_0.address
			WATCHDOG_TIMER_HW_IP_0_avalon_slave_0_write                => mm_interconnect_0_watchdog_timer_hw_ip_0_avalon_slave_0_write,      --                                                     .write
			WATCHDOG_TIMER_HW_IP_0_avalon_slave_0_read                 => mm_interconnect_0_watchdog_timer_hw_ip_0_avalon_slave_0_read,       --                                                     .read
			WATCHDOG_TIMER_HW_IP_0_avalon_slave_0_readdata             => mm_interconnect_0_watchdog_timer_hw_ip_0_avalon_slave_0_readdata,   --                                                     .readdata
			WATCHDOG_TIMER_HW_IP_0_avalon_slave_0_writedata            => mm_interconnect_0_watchdog_timer_hw_ip_0_avalon_slave_0_writedata,  --                                                     .writedata
			WATCHDOG_TIMER_HW_IP_0_avalon_slave_0_chipselect           => mm_interconnect_0_watchdog_timer_hw_ip_0_avalon_slave_0_chipselect  --                                                     .chipselect
		);

	irq_mapper : component watchdog_cpu_sys_irq_mapper
		port map (
			clk           => altpll_0_c0_clk,                --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			sender_irq    => cpu_irq_irq                     --    sender.irq
		);

	rst_controller : component watchdog_cpu_sys_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => cpu_debug_reset_request_reset,      -- reset_in1.reset
			clk            => altpll_0_c0_clk,                    --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_001 : component watchdog_cpu_sys_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => cpu_debug_reset_request_reset,      -- reset_in1.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;

	mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_chipselect_ports_inv <= not mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_chipselect;

	mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_read_ports_inv <= not mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_read;

	mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_write_ports_inv <= not mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_write;

	mm_interconnect_0_watchdog_timer_hw_ip_0_avalon_slave_0_chipselect_ports_inv <= not mm_interconnect_0_watchdog_timer_hw_ip_0_avalon_slave_0_chipselect;

	mm_interconnect_0_watchdog_timer_hw_ip_0_avalon_slave_0_read_ports_inv <= not mm_interconnect_0_watchdog_timer_hw_ip_0_avalon_slave_0_read;

	mm_interconnect_0_watchdog_timer_hw_ip_0_avalon_slave_0_write_ports_inv <= not mm_interconnect_0_watchdog_timer_hw_ip_0_avalon_slave_0_write;

	mm_interconnect_0_ledr_s1_write_ports_inv <= not mm_interconnect_0_ledr_s1_write;

	mm_interconnect_0_seven_seg_s1_write_ports_inv <= not mm_interconnect_0_seven_seg_s1_write;

	mm_interconnect_0_sdram_controller_s1_read_ports_inv <= not mm_interconnect_0_sdram_controller_s1_read;

	mm_interconnect_0_sdram_controller_s1_byteenable_ports_inv <= not mm_interconnect_0_sdram_controller_s1_byteenable;

	mm_interconnect_0_sdram_controller_s1_write_ports_inv <= not mm_interconnect_0_sdram_controller_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of watchdog_cpu_sys
