// ultrasonic_vga_system.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module ultrasonic_vga_system (
		input  wire        clk_clk,       //       clk.clk
		input  wire        reset_reset_n, //     reset.reset_n
		output wire [12:0] sdram_addr,    //     sdram.addr
		output wire [1:0]  sdram_ba,      //          .ba
		output wire        sdram_cas_n,   //          .cas_n
		output wire        sdram_cke,     //          .cke
		output wire        sdram_cs_n,    //          .cs_n
		inout  wire [15:0] sdram_dq,      //          .dq
		output wire [1:0]  sdram_dqm,     //          .dqm
		output wire        sdram_ras_n,   //          .ras_n
		output wire        sdram_we_n,    //          .we_n
		output wire        sdram_clk_clk, // sdram_clk.clk
		output wire [3:0]  vga_b_vga_b,   //     vga_b.vga_b
		output wire [3:0]  vga_g_vga_g,   //     vga_g.vga_g
		output wire        vga_hs_vga_hs, //    vga_hs.vga_hs
		output wire [3:0]  vga_r_vga_r,   //     vga_r.vga_r
		output wire        vga_vs_vga_vs  //    vga_vs.vga_vs
	);

	wire         altpll_0_c0_clk;                                         // altpll_0:c0 -> [VGA_IP_0:clk, irq_mapper:clk, jtag:clk, mm_interconnect_0:altpll_0_c0_clk, nios2_cpu:clk, rst_controller_002:clk, sdram_controller:clk, sram:clk, sysid_qsys_0:clock]
	wire         altpll_0_c2_clk;                                         // altpll_0:c2 -> [VGA_IP_0:clock_25, rst_controller:clk]
	wire  [31:0] nios2_cpu_data_master_readdata;                          // mm_interconnect_0:nios2_cpu_data_master_readdata -> nios2_cpu:d_readdata
	wire         nios2_cpu_data_master_waitrequest;                       // mm_interconnect_0:nios2_cpu_data_master_waitrequest -> nios2_cpu:d_waitrequest
	wire         nios2_cpu_data_master_debugaccess;                       // nios2_cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_cpu_data_master_debugaccess
	wire  [27:0] nios2_cpu_data_master_address;                           // nios2_cpu:d_address -> mm_interconnect_0:nios2_cpu_data_master_address
	wire   [3:0] nios2_cpu_data_master_byteenable;                        // nios2_cpu:d_byteenable -> mm_interconnect_0:nios2_cpu_data_master_byteenable
	wire         nios2_cpu_data_master_read;                              // nios2_cpu:d_read -> mm_interconnect_0:nios2_cpu_data_master_read
	wire         nios2_cpu_data_master_write;                             // nios2_cpu:d_write -> mm_interconnect_0:nios2_cpu_data_master_write
	wire  [31:0] nios2_cpu_data_master_writedata;                         // nios2_cpu:d_writedata -> mm_interconnect_0:nios2_cpu_data_master_writedata
	wire  [31:0] nios2_cpu_instruction_master_readdata;                   // mm_interconnect_0:nios2_cpu_instruction_master_readdata -> nios2_cpu:i_readdata
	wire         nios2_cpu_instruction_master_waitrequest;                // mm_interconnect_0:nios2_cpu_instruction_master_waitrequest -> nios2_cpu:i_waitrequest
	wire  [27:0] nios2_cpu_instruction_master_address;                    // nios2_cpu:i_address -> mm_interconnect_0:nios2_cpu_instruction_master_address
	wire         nios2_cpu_instruction_master_read;                       // nios2_cpu:i_read -> mm_interconnect_0:nios2_cpu_instruction_master_read
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_chipselect;     // mm_interconnect_0:jtag_avalon_jtag_slave_chipselect -> jtag:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_readdata;       // jtag:av_readdata -> mm_interconnect_0:jtag_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest;    // jtag:av_waitrequest -> mm_interconnect_0:jtag_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_avalon_jtag_slave_address;        // mm_interconnect_0:jtag_avalon_jtag_slave_address -> jtag:av_address
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_read;           // mm_interconnect_0:jtag_avalon_jtag_slave_read -> jtag:av_read_n
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_write;          // mm_interconnect_0:jtag_avalon_jtag_slave_write -> jtag:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_writedata;      // mm_interconnect_0:jtag_avalon_jtag_slave_writedata -> jtag:av_writedata
	wire         mm_interconnect_0_vga_ip_0_avalon_slave_0_chipselect;    // mm_interconnect_0:VGA_IP_0_avalon_slave_0_chipselect -> VGA_IP_0:cs_n
	wire  [31:0] mm_interconnect_0_vga_ip_0_avalon_slave_0_readdata;      // VGA_IP_0:dout -> mm_interconnect_0:VGA_IP_0_avalon_slave_0_readdata
	wire  [16:0] mm_interconnect_0_vga_ip_0_avalon_slave_0_address;       // mm_interconnect_0:VGA_IP_0_avalon_slave_0_address -> VGA_IP_0:addr
	wire         mm_interconnect_0_vga_ip_0_avalon_slave_0_read;          // mm_interconnect_0:VGA_IP_0_avalon_slave_0_read -> VGA_IP_0:read_n
	wire         mm_interconnect_0_vga_ip_0_avalon_slave_0_write;         // mm_interconnect_0:VGA_IP_0_avalon_slave_0_write -> VGA_IP_0:write_n
	wire  [31:0] mm_interconnect_0_vga_ip_0_avalon_slave_0_writedata;     // mm_interconnect_0:VGA_IP_0_avalon_slave_0_writedata -> VGA_IP_0:din
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;   // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;    // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire  [31:0] mm_interconnect_0_nios2_cpu_debug_mem_slave_readdata;    // nios2_cpu:debug_mem_slave_readdata -> mm_interconnect_0:nios2_cpu_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_cpu_debug_mem_slave_waitrequest; // nios2_cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_cpu_debug_mem_slave_debugaccess; // mm_interconnect_0:nios2_cpu_debug_mem_slave_debugaccess -> nios2_cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_cpu_debug_mem_slave_address;     // mm_interconnect_0:nios2_cpu_debug_mem_slave_address -> nios2_cpu:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_cpu_debug_mem_slave_read;        // mm_interconnect_0:nios2_cpu_debug_mem_slave_read -> nios2_cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_cpu_debug_mem_slave_byteenable;  // mm_interconnect_0:nios2_cpu_debug_mem_slave_byteenable -> nios2_cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_cpu_debug_mem_slave_write;       // mm_interconnect_0:nios2_cpu_debug_mem_slave_write -> nios2_cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_cpu_debug_mem_slave_writedata;   // mm_interconnect_0:nios2_cpu_debug_mem_slave_writedata -> nios2_cpu:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_altpll_0_pll_slave_readdata;           // altpll_0:readdata -> mm_interconnect_0:altpll_0_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_altpll_0_pll_slave_address;            // mm_interconnect_0:altpll_0_pll_slave_address -> altpll_0:address
	wire         mm_interconnect_0_altpll_0_pll_slave_read;               // mm_interconnect_0:altpll_0_pll_slave_read -> altpll_0:read
	wire         mm_interconnect_0_altpll_0_pll_slave_write;              // mm_interconnect_0:altpll_0_pll_slave_write -> altpll_0:write
	wire  [31:0] mm_interconnect_0_altpll_0_pll_slave_writedata;          // mm_interconnect_0:altpll_0_pll_slave_writedata -> altpll_0:writedata
	wire         mm_interconnect_0_sram_s1_chipselect;                    // mm_interconnect_0:sram_s1_chipselect -> sram:chipselect
	wire  [31:0] mm_interconnect_0_sram_s1_readdata;                      // sram:readdata -> mm_interconnect_0:sram_s1_readdata
	wire  [14:0] mm_interconnect_0_sram_s1_address;                       // mm_interconnect_0:sram_s1_address -> sram:address
	wire   [3:0] mm_interconnect_0_sram_s1_byteenable;                    // mm_interconnect_0:sram_s1_byteenable -> sram:byteenable
	wire         mm_interconnect_0_sram_s1_write;                         // mm_interconnect_0:sram_s1_write -> sram:write
	wire  [31:0] mm_interconnect_0_sram_s1_writedata;                     // mm_interconnect_0:sram_s1_writedata -> sram:writedata
	wire         mm_interconnect_0_sram_s1_clken;                         // mm_interconnect_0:sram_s1_clken -> sram:clken
	wire         mm_interconnect_0_sdram_controller_s1_chipselect;        // mm_interconnect_0:sdram_controller_s1_chipselect -> sdram_controller:az_cs
	wire  [15:0] mm_interconnect_0_sdram_controller_s1_readdata;          // sdram_controller:za_data -> mm_interconnect_0:sdram_controller_s1_readdata
	wire         mm_interconnect_0_sdram_controller_s1_waitrequest;       // sdram_controller:za_waitrequest -> mm_interconnect_0:sdram_controller_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_controller_s1_address;           // mm_interconnect_0:sdram_controller_s1_address -> sdram_controller:az_addr
	wire         mm_interconnect_0_sdram_controller_s1_read;              // mm_interconnect_0:sdram_controller_s1_read -> sdram_controller:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_controller_s1_byteenable;        // mm_interconnect_0:sdram_controller_s1_byteenable -> sdram_controller:az_be_n
	wire         mm_interconnect_0_sdram_controller_s1_readdatavalid;     // sdram_controller:za_valid -> mm_interconnect_0:sdram_controller_s1_readdatavalid
	wire         mm_interconnect_0_sdram_controller_s1_write;             // mm_interconnect_0:sdram_controller_s1_write -> sdram_controller:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_controller_s1_writedata;         // mm_interconnect_0:sdram_controller_s1_writedata -> sdram_controller:az_data
	wire         irq_mapper_receiver0_irq;                                // jtag:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2_cpu_irq_irq;                                       // irq_mapper:sender_irq -> nios2_cpu:irq
	wire         rst_controller_reset_out_reset;                          // rst_controller:reset_out -> VGA_IP_0:reset_n
	wire         nios2_cpu_debug_reset_request_reset;                     // nios2_cpu:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_002:reset_in1]
	wire         rst_controller_001_reset_out_reset;                      // rst_controller_001:reset_out -> [altpll_0:reset, mm_interconnect_0:altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_002_reset_out_reset;                      // rst_controller_002:reset_out -> [irq_mapper:reset, jtag:rst_n, mm_interconnect_0:nios2_cpu_reset_reset_bridge_in_reset_reset, nios2_cpu:reset_n, rst_translator:in_reset, sdram_controller:reset_n, sram:reset, sysid_qsys_0:reset_n]
	wire         rst_controller_002_reset_out_reset_req;                  // rst_controller_002:reset_req -> [nios2_cpu:reset_req, rst_translator:reset_req_in, sram:reset_req]

	VGA_IP vga_ip_0 (
		.clk      (altpll_0_c0_clk),                                       //          clock.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //          reset.reset_n
		.addr     (mm_interconnect_0_vga_ip_0_avalon_slave_0_address),     // avalon_slave_0.address
		.cs_n     (~mm_interconnect_0_vga_ip_0_avalon_slave_0_chipselect), //               .chipselect_n
		.read_n   (~mm_interconnect_0_vga_ip_0_avalon_slave_0_read),       //               .read_n
		.write_n  (~mm_interconnect_0_vga_ip_0_avalon_slave_0_write),      //               .write_n
		.din      (mm_interconnect_0_vga_ip_0_avalon_slave_0_writedata),   //               .writedata
		.dout     (mm_interconnect_0_vga_ip_0_avalon_slave_0_readdata),    //               .readdata
		.clock_25 (altpll_0_c2_clk),                                       //  clock_sink_25.clk
		.vga_b    (vga_b_vga_b),                                           //  conduit_end_1.vga_b
		.vga_g    (vga_g_vga_g),                                           //  conduit_end_2.vga_g
		.vga_hs   (vga_hs_vga_hs),                                         //  conduit_end_3.vga_hs
		.vga_r    (vga_r_vga_r),                                           //  conduit_end_4.vga_r
		.vga_vs   (vga_vs_vga_vs)                                          //  conduit_end_5.vga_vs
	);

	ultrasonic_vga_system_altpll_0 altpll_0 (
		.clk                (clk_clk),                                        //       inclk_interface.clk
		.reset              (rst_controller_001_reset_out_reset),             // inclk_interface_reset.reset
		.read               (mm_interconnect_0_altpll_0_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_altpll_0_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_altpll_0_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_altpll_0_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_altpll_0_pll_slave_writedata), //                      .writedata
		.c0                 (altpll_0_c0_clk),                                //                    c0.clk
		.c1                 (sdram_clk_clk),                                  //                    c1.clk
		.c2                 (altpll_0_c2_clk),                                //                    c2.clk
		.scandone           (),                                               //           (terminated)
		.scandataout        (),                                               //           (terminated)
		.c3                 (),                                               //           (terminated)
		.c4                 (),                                               //           (terminated)
		.areset             (1'b0),                                           //           (terminated)
		.locked             (),                                               //           (terminated)
		.phasedone          (),                                               //           (terminated)
		.phasecounterselect (3'b000),                                         //           (terminated)
		.phaseupdown        (1'b0),                                           //           (terminated)
		.phasestep          (1'b0),                                           //           (terminated)
		.scanclk            (1'b0),                                           //           (terminated)
		.scanclkena         (1'b0),                                           //           (terminated)
		.scandata           (1'b0),                                           //           (terminated)
		.configupdate       (1'b0)                                            //           (terminated)
	);

	ultrasonic_vga_system_jtag jtag (
		.clk            (altpll_0_c0_clk),                                      //               clk.clk
		.rst_n          (~rst_controller_002_reset_out_reset),                  //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                              //               irq.irq
	);

	ultrasonic_vga_system_nios2_cpu nios2_cpu (
		.clk                                 (altpll_0_c0_clk),                                         //                       clk.clk
		.reset_n                             (~rst_controller_002_reset_out_reset),                     //                     reset.reset_n
		.reset_req                           (rst_controller_002_reset_out_reset_req),                  //                          .reset_req
		.d_address                           (nios2_cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_cpu_data_master_read),                              //                          .read
		.d_readdata                          (nios2_cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_cpu_data_master_write),                             //                          .write
		.d_writedata                         (nios2_cpu_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_cpu_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_cpu_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                         // custom_instruction_master.readra
	);

	ultrasonic_vga_system_sdram_controller sdram_controller (
		.clk            (altpll_0_c0_clk),                                     //   clk.clk
		.reset_n        (~rst_controller_002_reset_out_reset),                 // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_controller_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_controller_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_controller_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_controller_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_controller_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_controller_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_controller_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_controller_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_controller_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                                          //  wire.export
		.zs_ba          (sdram_ba),                                            //      .export
		.zs_cas_n       (sdram_cas_n),                                         //      .export
		.zs_cke         (sdram_cke),                                           //      .export
		.zs_cs_n        (sdram_cs_n),                                          //      .export
		.zs_dq          (sdram_dq),                                            //      .export
		.zs_dqm         (sdram_dqm),                                           //      .export
		.zs_ras_n       (sdram_ras_n),                                         //      .export
		.zs_we_n        (sdram_we_n)                                           //      .export
	);

	ultrasonic_vga_system_sram sram (
		.clk        (altpll_0_c0_clk),                        //   clk1.clk
		.address    (mm_interconnect_0_sram_s1_address),      //     s1.address
		.clken      (mm_interconnect_0_sram_s1_clken),        //       .clken
		.chipselect (mm_interconnect_0_sram_s1_chipselect),   //       .chipselect
		.write      (mm_interconnect_0_sram_s1_write),        //       .write
		.readdata   (mm_interconnect_0_sram_s1_readdata),     //       .readdata
		.writedata  (mm_interconnect_0_sram_s1_writedata),    //       .writedata
		.byteenable (mm_interconnect_0_sram_s1_byteenable),   //       .byteenable
		.reset      (rst_controller_002_reset_out_reset),     // reset1.reset
		.reset_req  (rst_controller_002_reset_out_reset_req), //       .reset_req
		.freeze     (1'b0)                                    // (terminated)
	);

	ultrasonic_vga_system_sysid_qsys_0 sysid_qsys_0 (
		.clock    (altpll_0_c0_clk),                                       //           clk.clk
		.reset_n  (~rst_controller_002_reset_out_reset),                   //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	ultrasonic_vga_system_mm_interconnect_0 mm_interconnect_0 (
		.altpll_0_c0_clk                                            (altpll_0_c0_clk),                                         //                                          altpll_0_c0.clk
		.clk_0_clk_clk                                              (clk_clk),                                                 //                                            clk_0_clk.clk
		.altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                      // altpll_0_inclk_interface_reset_reset_bridge_in_reset.reset
		.nios2_cpu_reset_reset_bridge_in_reset_reset                (rst_controller_002_reset_out_reset),                      //                nios2_cpu_reset_reset_bridge_in_reset.reset
		.nios2_cpu_data_master_address                              (nios2_cpu_data_master_address),                           //                                nios2_cpu_data_master.address
		.nios2_cpu_data_master_waitrequest                          (nios2_cpu_data_master_waitrequest),                       //                                                     .waitrequest
		.nios2_cpu_data_master_byteenable                           (nios2_cpu_data_master_byteenable),                        //                                                     .byteenable
		.nios2_cpu_data_master_read                                 (nios2_cpu_data_master_read),                              //                                                     .read
		.nios2_cpu_data_master_readdata                             (nios2_cpu_data_master_readdata),                          //                                                     .readdata
		.nios2_cpu_data_master_write                                (nios2_cpu_data_master_write),                             //                                                     .write
		.nios2_cpu_data_master_writedata                            (nios2_cpu_data_master_writedata),                         //                                                     .writedata
		.nios2_cpu_data_master_debugaccess                          (nios2_cpu_data_master_debugaccess),                       //                                                     .debugaccess
		.nios2_cpu_instruction_master_address                       (nios2_cpu_instruction_master_address),                    //                         nios2_cpu_instruction_master.address
		.nios2_cpu_instruction_master_waitrequest                   (nios2_cpu_instruction_master_waitrequest),                //                                                     .waitrequest
		.nios2_cpu_instruction_master_read                          (nios2_cpu_instruction_master_read),                       //                                                     .read
		.nios2_cpu_instruction_master_readdata                      (nios2_cpu_instruction_master_readdata),                   //                                                     .readdata
		.altpll_0_pll_slave_address                                 (mm_interconnect_0_altpll_0_pll_slave_address),            //                                   altpll_0_pll_slave.address
		.altpll_0_pll_slave_write                                   (mm_interconnect_0_altpll_0_pll_slave_write),              //                                                     .write
		.altpll_0_pll_slave_read                                    (mm_interconnect_0_altpll_0_pll_slave_read),               //                                                     .read
		.altpll_0_pll_slave_readdata                                (mm_interconnect_0_altpll_0_pll_slave_readdata),           //                                                     .readdata
		.altpll_0_pll_slave_writedata                               (mm_interconnect_0_altpll_0_pll_slave_writedata),          //                                                     .writedata
		.jtag_avalon_jtag_slave_address                             (mm_interconnect_0_jtag_avalon_jtag_slave_address),        //                               jtag_avalon_jtag_slave.address
		.jtag_avalon_jtag_slave_write                               (mm_interconnect_0_jtag_avalon_jtag_slave_write),          //                                                     .write
		.jtag_avalon_jtag_slave_read                                (mm_interconnect_0_jtag_avalon_jtag_slave_read),           //                                                     .read
		.jtag_avalon_jtag_slave_readdata                            (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),       //                                                     .readdata
		.jtag_avalon_jtag_slave_writedata                           (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),      //                                                     .writedata
		.jtag_avalon_jtag_slave_waitrequest                         (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest),    //                                                     .waitrequest
		.jtag_avalon_jtag_slave_chipselect                          (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),     //                                                     .chipselect
		.nios2_cpu_debug_mem_slave_address                          (mm_interconnect_0_nios2_cpu_debug_mem_slave_address),     //                            nios2_cpu_debug_mem_slave.address
		.nios2_cpu_debug_mem_slave_write                            (mm_interconnect_0_nios2_cpu_debug_mem_slave_write),       //                                                     .write
		.nios2_cpu_debug_mem_slave_read                             (mm_interconnect_0_nios2_cpu_debug_mem_slave_read),        //                                                     .read
		.nios2_cpu_debug_mem_slave_readdata                         (mm_interconnect_0_nios2_cpu_debug_mem_slave_readdata),    //                                                     .readdata
		.nios2_cpu_debug_mem_slave_writedata                        (mm_interconnect_0_nios2_cpu_debug_mem_slave_writedata),   //                                                     .writedata
		.nios2_cpu_debug_mem_slave_byteenable                       (mm_interconnect_0_nios2_cpu_debug_mem_slave_byteenable),  //                                                     .byteenable
		.nios2_cpu_debug_mem_slave_waitrequest                      (mm_interconnect_0_nios2_cpu_debug_mem_slave_waitrequest), //                                                     .waitrequest
		.nios2_cpu_debug_mem_slave_debugaccess                      (mm_interconnect_0_nios2_cpu_debug_mem_slave_debugaccess), //                                                     .debugaccess
		.sdram_controller_s1_address                                (mm_interconnect_0_sdram_controller_s1_address),           //                                  sdram_controller_s1.address
		.sdram_controller_s1_write                                  (mm_interconnect_0_sdram_controller_s1_write),             //                                                     .write
		.sdram_controller_s1_read                                   (mm_interconnect_0_sdram_controller_s1_read),              //                                                     .read
		.sdram_controller_s1_readdata                               (mm_interconnect_0_sdram_controller_s1_readdata),          //                                                     .readdata
		.sdram_controller_s1_writedata                              (mm_interconnect_0_sdram_controller_s1_writedata),         //                                                     .writedata
		.sdram_controller_s1_byteenable                             (mm_interconnect_0_sdram_controller_s1_byteenable),        //                                                     .byteenable
		.sdram_controller_s1_readdatavalid                          (mm_interconnect_0_sdram_controller_s1_readdatavalid),     //                                                     .readdatavalid
		.sdram_controller_s1_waitrequest                            (mm_interconnect_0_sdram_controller_s1_waitrequest),       //                                                     .waitrequest
		.sdram_controller_s1_chipselect                             (mm_interconnect_0_sdram_controller_s1_chipselect),        //                                                     .chipselect
		.sram_s1_address                                            (mm_interconnect_0_sram_s1_address),                       //                                              sram_s1.address
		.sram_s1_write                                              (mm_interconnect_0_sram_s1_write),                         //                                                     .write
		.sram_s1_readdata                                           (mm_interconnect_0_sram_s1_readdata),                      //                                                     .readdata
		.sram_s1_writedata                                          (mm_interconnect_0_sram_s1_writedata),                     //                                                     .writedata
		.sram_s1_byteenable                                         (mm_interconnect_0_sram_s1_byteenable),                    //                                                     .byteenable
		.sram_s1_chipselect                                         (mm_interconnect_0_sram_s1_chipselect),                    //                                                     .chipselect
		.sram_s1_clken                                              (mm_interconnect_0_sram_s1_clken),                         //                                                     .clken
		.sysid_qsys_0_control_slave_address                         (mm_interconnect_0_sysid_qsys_0_control_slave_address),    //                           sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata                        (mm_interconnect_0_sysid_qsys_0_control_slave_readdata),   //                                                     .readdata
		.VGA_IP_0_avalon_slave_0_address                            (mm_interconnect_0_vga_ip_0_avalon_slave_0_address),       //                              VGA_IP_0_avalon_slave_0.address
		.VGA_IP_0_avalon_slave_0_write                              (mm_interconnect_0_vga_ip_0_avalon_slave_0_write),         //                                                     .write
		.VGA_IP_0_avalon_slave_0_read                               (mm_interconnect_0_vga_ip_0_avalon_slave_0_read),          //                                                     .read
		.VGA_IP_0_avalon_slave_0_readdata                           (mm_interconnect_0_vga_ip_0_avalon_slave_0_readdata),      //                                                     .readdata
		.VGA_IP_0_avalon_slave_0_writedata                          (mm_interconnect_0_vga_ip_0_avalon_slave_0_writedata),     //                                                     .writedata
		.VGA_IP_0_avalon_slave_0_chipselect                         (mm_interconnect_0_vga_ip_0_avalon_slave_0_chipselect)     //                                                     .chipselect
	);

	ultrasonic_vga_system_irq_mapper irq_mapper (
		.clk           (altpll_0_c0_clk),                    //       clk.clk
		.reset         (rst_controller_002_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.sender_irq    (nios2_cpu_irq_irq)                   //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                      // reset_in0.reset
		.reset_in1      (nios2_cpu_debug_reset_request_reset), // reset_in1.reset
		.clk            (altpll_0_c2_clk),                     //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),      // reset_out.reset
		.reset_req      (),                                    // (terminated)
		.reset_req_in0  (1'b0),                                // (terminated)
		.reset_req_in1  (1'b0),                                // (terminated)
		.reset_in2      (1'b0),                                // (terminated)
		.reset_req_in2  (1'b0),                                // (terminated)
		.reset_in3      (1'b0),                                // (terminated)
		.reset_req_in3  (1'b0),                                // (terminated)
		.reset_in4      (1'b0),                                // (terminated)
		.reset_req_in4  (1'b0),                                // (terminated)
		.reset_in5      (1'b0),                                // (terminated)
		.reset_req_in5  (1'b0),                                // (terminated)
		.reset_in6      (1'b0),                                // (terminated)
		.reset_req_in6  (1'b0),                                // (terminated)
		.reset_in7      (1'b0),                                // (terminated)
		.reset_req_in7  (1'b0),                                // (terminated)
		.reset_in8      (1'b0),                                // (terminated)
		.reset_req_in8  (1'b0),                                // (terminated)
		.reset_in9      (1'b0),                                // (terminated)
		.reset_req_in9  (1'b0),                                // (terminated)
		.reset_in10     (1'b0),                                // (terminated)
		.reset_req_in10 (1'b0),                                // (terminated)
		.reset_in11     (1'b0),                                // (terminated)
		.reset_req_in11 (1'b0),                                // (terminated)
		.reset_in12     (1'b0),                                // (terminated)
		.reset_req_in12 (1'b0),                                // (terminated)
		.reset_in13     (1'b0),                                // (terminated)
		.reset_req_in13 (1'b0),                                // (terminated)
		.reset_in14     (1'b0),                                // (terminated)
		.reset_req_in14 (1'b0),                                // (terminated)
		.reset_in15     (1'b0),                                // (terminated)
		.reset_req_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                      // reset_in0.reset
		.reset_in1      (nios2_cpu_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                             //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),  // reset_out.reset
		.reset_req      (),                                    // (terminated)
		.reset_req_in0  (1'b0),                                // (terminated)
		.reset_req_in1  (1'b0),                                // (terminated)
		.reset_in2      (1'b0),                                // (terminated)
		.reset_req_in2  (1'b0),                                // (terminated)
		.reset_in3      (1'b0),                                // (terminated)
		.reset_req_in3  (1'b0),                                // (terminated)
		.reset_in4      (1'b0),                                // (terminated)
		.reset_req_in4  (1'b0),                                // (terminated)
		.reset_in5      (1'b0),                                // (terminated)
		.reset_req_in5  (1'b0),                                // (terminated)
		.reset_in6      (1'b0),                                // (terminated)
		.reset_req_in6  (1'b0),                                // (terminated)
		.reset_in7      (1'b0),                                // (terminated)
		.reset_req_in7  (1'b0),                                // (terminated)
		.reset_in8      (1'b0),                                // (terminated)
		.reset_req_in8  (1'b0),                                // (terminated)
		.reset_in9      (1'b0),                                // (terminated)
		.reset_req_in9  (1'b0),                                // (terminated)
		.reset_in10     (1'b0),                                // (terminated)
		.reset_req_in10 (1'b0),                                // (terminated)
		.reset_in11     (1'b0),                                // (terminated)
		.reset_req_in11 (1'b0),                                // (terminated)
		.reset_in12     (1'b0),                                // (terminated)
		.reset_req_in12 (1'b0),                                // (terminated)
		.reset_in13     (1'b0),                                // (terminated)
		.reset_req_in13 (1'b0),                                // (terminated)
		.reset_in14     (1'b0),                                // (terminated)
		.reset_req_in14 (1'b0),                                // (terminated)
		.reset_in15     (1'b0),                                // (terminated)
		.reset_req_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_cpu_debug_reset_request_reset),    // reset_in1.reset
		.clk            (altpll_0_c0_clk),                        //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_002_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
